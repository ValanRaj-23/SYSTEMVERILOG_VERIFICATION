package my_pkg;
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "score_board.sv"
parameter int t = 20;
endpackage
