interface intf(input bit clk);
  logic rst;
  logic d;
  logic q;
  
  modport ds(input clk, rst, d, output q);
  modport tb(input q, output  rst, d);
  
endinterface
