temp.sv
